`ifndef __HAZARD_SV
`define __HAZARD_SV

`ifdef VERILATOR
`include "include/common.sv"
`include "include/pipes.sv"
`endif

module hazard
    import common::*;
    import pipes::*;(
    
);
    
endmodule

`endif
